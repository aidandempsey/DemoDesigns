-- Package
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
package MainPackage is


end MainPackage;
package body MainPackage is
end MainPackage;
